.subckt CLK_COMP clk clkbo dn dp gt vb vdd vin vinb vintn<2> vintn<1> vintp<2> vintp<1> vss
xm103 clkb clk vdd vdd pfet_lvt w=480e-9 l=40e-9 nf=1
xm30 clk net030 vdd vdd pfet_lvt w=3.84e-6 l=40e-9 nf=8
xm124 clkbo clk vdd vdd pfet_lvt w=480e-9 l=40e-9 nf=1
xm16 v2p vxn vdd _net0 pfet_lvt w=2.88e-6 l=40e-9 nf=6
xm114 d v2n vdd vdd pfet_lvt w=1.92e-6 l=40e-9 nf=4
xm122 dp db vdd vdd pfet_lvt w=960e-9 l=40e-9 nf=2
xm25 vmid v2p vdd vdd pfet_lvt w=960e-9 l=40e-9 nf=2
xm14 net027 d vdd vdd pfet_lvt w=480e-9 l=40e-9 nf=1
xm24 db v2p vdd vdd pfet_lvt w=1.92e-6 l=40e-9 nf=4
xm85 net030 gt vdd vdd pfet_lvt w=1.92e-6 l=40e-9 nf=2
xm6 net031 net027 vdd vdd pfet_lvt w=960e-9 l=40e-9 nf=1
xm8 db d vdd vdd pfet_lvt w=1.92e-6 l=40e-9 nf=4
xm5 d db vdd vdd pfet_lvt w=1.92e-6 l=40e-9 nf=4
xm119 dn d vdd vdd pfet_lvt w=960e-9 l=40e-9 nf=2
xm71 net027 db vdd vdd pfet_lvt w=480e-9 l=40e-9 nf=1
xm9 net030 net031 vdd vdd pfet_lvt w=1.92e-6 l=40e-9 nf=2
xm35 vxn clk vdd vdd pfet_lvt w=2.88e-6 l=40e-9 nf=6
xm73 vxp clk vdd vdd pfet_lvt w=2.88e-6 l=40e-9 nf=6
xm19 v2n vxp vdd _net0 pfet_lvt w=2.88e-6 l=40e-9 nf=6
xm26 vmidb v2n vdd vdd pfet_lvt w=960e-9 l=40e-9 nf=2
xm10 net030 net031 net032 vss nfet_lvt w=1.92e-6 l=40e-9 nf=4
xm69 v1p vintn<1> vss vss nfet_lvt w=720e-9 l=40e-9 nf=3
xm17 net032 gt vss vss nfet_lvt w=1.92e-6 l=40e-9 nf=4
xm116 vxp clk v1p vss nfet_lvt w=1.92e-6 l=40e-9 nf=4
xm102 clkb clk vss vss nfet_lvt w=240e-9 l=40e-9 nf=1
xm120 dn d vss vss nfet_lvt w=480e-9 l=40e-9 nf=1
xm1 db d vmid vss nfet_lvt w=1.92e-6 l=40e-9 nf=4
xm113 vmidb v2n vss vss nfet_lvt w=1.92e-6 l=40e-9 nf=4
xm7 net031 net027 vss vss nfet_lvt w=480e-9 l=40e-9 nf=1
xm28 vss vss v1p vss nfet_lvt w=240e-9 l=40e-9 nf=1
xm70 v1p vinb vss vss nfet_lvt w=240e-9 l=40e-9 nf=1
xm97 net027 clkb net0107 vss nfet_lvt w=480e-9 l=40e-9 nf=1
xm12 net0107 vb vss vss nfet_lvt w=1.92e-6 l=40e-9 nf=4
xm121 dp db vss vss nfet_lvt w=480e-9 l=40e-9 nf=1
xm115 vxn clk v1n vss nfet_lvt w=1.92e-6 l=40e-9 nf=4
xm27 clk net030 vss vss nfet_lvt w=1.92e-6 l=40e-9 nf=2
xm20 v2p vxn vss vss nfet_lvt w=1.92e-6 l=40e-9 nf=4
xm3 d db vmidb vss nfet_lvt w=1.92e-6 l=40e-9 nf=4
xm18 vss vss vss vss nfet_lvt w=240e-9 l=40e-9 nf=1
xm55 v1n vin vss vss nfet_lvt w=240e-9 l=40e-9 nf=1
xm23 vss vss v1n vss nfet_lvt w=240e-9 l=40e-9 nf=1
xm57 v1n vintp<2> vss vss nfet_lvt w=2.88e-6 l=40e-9 nf=12
xm125 clkbo clk vss vss nfet_lvt w=240e-9 l=40e-9 nf=1
xm22 vmid v2p vss vss nfet_lvt w=1.92e-6 l=40e-9 nf=4
xm21 v2n vxp vss vss nfet_lvt w=1.92e-6 l=40e-9 nf=4
xm56 v1n vintp<1> vss vss nfet_lvt w=720e-9 l=40e-9 nf=3
xm68 v1p vintn<2> vss vss nfet_lvt w=2.88e-6 l=40e-9 nf=12
.ends CLK_COMP
