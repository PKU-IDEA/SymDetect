.subckt C1 a b vss
xc0<3> a b vss cap
xc0<2> a b vss cap
xc0<1> a b vss cap
xc0<0> a b vss cap
.ends C1